module invert(input signal, output out);
  assign out = ~signal;
endmodule
